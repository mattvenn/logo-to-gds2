VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LOGO
  CLASS block ;
  FOREIGN LOGO ;
  ORIGIN -462.900 1677.010 ;
  SIZE 390.420 BY 280.970 ;
  SYMMETRY X Y R90 ;
  OBS
      LAYER met4 ;
        RECT 540.000 -1462.560 555.000 -1453.560 ;
        RECT 591.000 -1462.560 606.000 -1453.560 ;
        RECT 540.000 -1483.560 606.000 -1462.560 ;
        RECT 540.000 -1530.000 555.000 -1483.560 ;
        RECT 567.000 -1498.560 579.000 -1483.560 ;
        RECT 591.000 -1530.000 606.000 -1483.560 ;
        RECT 618.000 -1470.000 663.000 -1453.560 ;
        RECT 675.000 -1470.000 720.000 -1455.000 ;
        RECT 735.000 -1470.000 780.000 -1455.000 ;
        RECT 618.000 -1485.000 633.000 -1470.000 ;
        RECT 648.000 -1485.000 663.000 -1470.000 ;
        RECT 618.000 -1500.000 663.000 -1485.000 ;
        RECT 618.000 -1530.000 633.000 -1500.000 ;
        RECT 648.000 -1530.000 663.000 -1500.000 ;
        RECT 690.000 -1530.000 705.000 -1470.000 ;
        RECT 750.000 -1530.000 765.000 -1470.000 ;
        RECT 540.000 -1597.560 555.000 -1545.000 ;
        RECT 591.000 -1597.560 606.000 -1545.000 ;
        RECT 540.000 -1618.560 606.000 -1597.560 ;
        RECT 615.000 -1560.000 660.000 -1545.000 ;
        RECT 615.000 -1575.000 630.000 -1560.000 ;
        RECT 669.000 -1561.560 684.000 -1546.560 ;
        RECT 705.000 -1561.560 720.000 -1546.560 ;
        RECT 669.000 -1573.560 720.000 -1561.560 ;
        RECT 615.000 -1590.000 645.000 -1575.000 ;
        RECT 615.000 -1605.000 630.000 -1590.000 ;
        RECT 615.000 -1618.560 660.000 -1605.000 ;
        RECT 669.000 -1618.560 684.000 -1573.560 ;
        RECT 705.000 -1618.560 720.000 -1573.560 ;
        RECT 729.000 -1561.560 744.000 -1546.560 ;
        RECT 765.000 -1561.560 780.000 -1546.560 ;
        RECT 729.000 -1573.560 780.000 -1561.560 ;
        RECT 729.000 -1618.560 744.000 -1573.560 ;
        RECT 765.000 -1618.560 780.000 -1573.560 ;
  END
END LOGO
END LIBRARY

