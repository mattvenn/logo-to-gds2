VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LOGO
  CLASS BLOCK ;
  FOREIGN LOGO ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.005 BY 0.005 ;
END LOGO
END LIBRARY

